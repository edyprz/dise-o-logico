--Edgar Humberto Perez Martinez
--Ing Electronica
--Descripcion de un decodificador bcd de 7 segmentos  
entity decobcd7seg is
   port( 

	ent: in bit_vector(3 downto 0);
	sal: out bit_vector(6 downto 0)
       );
end entity decobcd7seg;

architecture beh of decobcd7seg is
begin

   sal <= "1111110" when ent = "0000" else
	  "0110000" when ent = "0001" else
	  "1101101" when ent = "0010" else
	  "1111001" when ent = "0011" else
	  "0110011" when ent = "0100" else
          "1011011" when ent = "0101" else
          "1011111" when ent = "0110" else
	  "1110000" when ent = "0111" else
          "1111111" when ent = "1000" else
          "1111011" when ent = "1001" else
          "1001111" ;


end architecture beh;
				
